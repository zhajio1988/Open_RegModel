`define PICO_FEATURE_DATA_TYPE_INT8
`define PICO_BPE 8
`define PICO_WEIGHT_DATA_TYPE_INT8
`define PICO_SDP_BS_ENABLE
`define PICO_SDP_BN_ENABLE
`define PICO_PDP_ENABLE
`define PICO_CDP_ENABLE
`define PICO_MAC_ATOMIC_C_SIZE 32
`define PICO_MAC_ATOMIC_K_SIZE 8
`define PICO_MEMORY_ATOMIC_SIZE 8
`define PICO_CBUF_BANK_NUMBER 32
`define PICO_CBUF_BANK_WIDTH 32
`define PICO_CBUF_BANK_DEPTH 128
`define PICO_SDP_BS_THROUGHPUT 1
`define PICO_SDP_BN_THROUGHPUT 1
`define PICO_SDP_EW_THROUGHPUT 0
`define PICO_SDP_EW_THROUGHPUT_LOG2 0
`define PICO_SDP_MAX_THROUGHPUT 1
`define PICO_SDP2PDP_WIDTH 8
`define PICO_PDP_THROUGHPUT 1
`define PICO_CDP_THROUGHPUT 1
`define PICO_PRIMARY_MEMIF_LATENCY 64
`define PICO_PRIMARY_MEMIF_MAX_BURST_LENGTH 1
`define PICO_PRIMARY_MEMIF_WIDTH 64
`define PICO_MEM_ADDRESS_WIDTH 32
`define PICO_MEMIF_WIDTH 64
`define PICO_DMA_RD_SIZE 15
`define PICO_DMA_WR_SIZE 13
`define PICO_DMA_MASK_BIT 1
`define PICO_DMA_RD_RSP 65
`define PICO_DMA_WR_REQ 66
`define PICO_DMA_WR_CMD 46
`define PICO_DMA_RD_REQ 47
`define PICO_MEMORY_ATOMIC_LOG2 3
`define PICO_PRIMARY_MEMIF_WIDTH_LOG2 3
`define PICO_MEMORY_ATOMIC_WIDTH 64
`define PICO_MCIF_BURST_SIZE 1
`define PICO_MCIF_BURST_SIZE_LOG2 0
`define PICO_NUM_DMA_READ_CLIENTS 7
`define PICO_NUM_DMA_WRITE_CLIENTS 3
`define PDP_SINGLE_LBUF_WIDTH 128
`define PDP_SINGLE_LBUF_DEPTH 14
`define PICO_VMOD_PRIMARY_BANDWIDTH 2
`define PICO_VMOD_SDP_MRDMA_OUTPUT_THROUGHPUT 1
`define PICO_VMOD_SDP_BRDMA_OUTPUT_THROUGHPUT 4
`define PICO_VMOD_SDP_NRDMA_OUTPUT_THROUGHPUT 4
`define PICO_VMOD_SDP_ERDMA_OUTPUT_THROUGHPUT 0
`define PICO_VMOD_CDP_RDMA_OUTPUT_THROUGHPUT_USE 1
`define PICO_VMOD_PDP_RDMA_OUTPUT_THROUGHPUT_USE 1
`define PICO_VMOD_SDP_MRDMA_OUTPUT_THROUGHPUT_USE 1
`define PICO_VMOD_SDP_BRDMA_OUTPUT_THROUGHPUT_USE 2
`define PICO_VMOD_SDP_NRDMA_OUTPUT_THROUGHPUT_USE 2
`define PICO_VMOD_SDP_ERDMA_OUTPUT_THROUGHPUT_USE 0
`define PICO_VMOD_CDP_RDMA_LATENCY_FIFO_DEPTH 8
`define PICO_VMOD_PDP_RDMA_LATENCY_FIFO_DEPTH 8
`define PICO_VMOD_SDP_MRDMA_LATENCY_FIFO_DEPTH 8
`define PICO_VMOD_SDP_BRDMA_LATENCY_FIFO_DEPTH 16
`define PICO_VMOD_SDP_NRDMA_LATENCY_FIFO_DEPTH 16
`define PICO_VMOD_SDP_ERDMA_LATENCY_FIFO_DEPTH 4
`define PICO_VMOD_DMA_LAT_FIFO_DEPTH_MAX 512
`define PICO_MAC_ATOMIC_C_SIZE_LOG2 5
`define PICO_MAC_ATOMIC_K_SIZE_LOG2 3
`define PICO_MAC_ATOMIC_K_SIZE_DIV2 4
`define PICO_CBUF_BANK_NUMBER_LOG2 5
`define PICO_CBUF_BANK_WIDTH_LOG2 5
`define PICO_CBUF_BANK_DEPTH_LOG2 7
`define PICO_CBUF_DEPTH_LOG2 12
`define PICO_CBUF_ENTRY_WIDTH 256
`define PICO_CBUF_WIDTH_LOG2 8
`define PICO_CBUF_WIDTH_MUL2_LOG2 9
`define PICO_BPE_LOG2 3
`define PICO_MAC_RESULT_WIDTH 21
`define PICO_CC_ATOMC_DIV_ATOMK 4
`define PICO_CACC_SDP_WIDTH 34
`define PICO_CACC_SDP_SINGLE_THROUGHPUT 32
`define PICO_CDMA_GRAIN_MAX_BIT 13